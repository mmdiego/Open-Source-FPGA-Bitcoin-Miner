
// Generate a clock to be used by the hashing cores.

module hashing_pll # (
	parameter INPUT_FREQUENCY = 50,
	parameter DIVIDE_BY = 1,
	parameter MULTIPLY_BY = 1
) (
	input areset,
	input rx_clk,
	output [1:0] tx_hash_clk,
	output lock
);

//	wire [4:0] clks;
//
//	assign tx_hash_clk = clks[0];

	altera_pll #(
		.fractional_vco_multiplier("false"),
		.reference_clock_frequency((1000000 / INPUT_FREQUENCY)),
		.operation_mode("direct"),
		.number_of_clocks(2),
		.output_clock_frequency0((1000000 * DIVIDE_BY) / (INPUT_FREQUENCY * MULTIPLY_BY)),
		.phase_shift0("0 ps"),
		.duty_cycle0(50),
		.output_clock_frequency1((1000000 * DIVIDE_BY) / (INPUT_FREQUENCY * 2 * MULTIPLY_BY)),
		.phase_shift1("0 ps"),
		.duty_cycle1(50),
		.output_clock_frequency2("0 MHz"),
		.phase_shift2("0 ps"),
		.duty_cycle2(50),
		.output_clock_frequency3("0 MHz"),
		.phase_shift3("0 ps"),
		.duty_cycle3(50),
		.output_clock_frequency4("0 MHz"),
		.phase_shift4("0 ps"),
		.duty_cycle4(50),
		.output_clock_frequency5("0 MHz"),
		.phase_shift5("0 ps"),
		.duty_cycle5(50),
		.output_clock_frequency6("0 MHz"),
		.phase_shift6("0 ps"),
		.duty_cycle6(50),
		.output_clock_frequency7("0 MHz"),
		.phase_shift7("0 ps"),
		.duty_cycle7(50),
		.output_clock_frequency8("0 MHz"),
		.phase_shift8("0 ps"),
		.duty_cycle8(50),
		.output_clock_frequency9("0 MHz"),
		.phase_shift9("0 ps"),
		.duty_cycle9(50),
		.output_clock_frequency10("0 MHz"),
		.phase_shift10("0 ps"),
		.duty_cycle10(50),
		.output_clock_frequency11("0 MHz"),
		.phase_shift11("0 ps"),
		.duty_cycle11(50),
		.output_clock_frequency12("0 MHz"),
		.phase_shift12("0 ps"),
		.duty_cycle12(50),
		.output_clock_frequency13("0 MHz"),
		.phase_shift13("0 ps"),
		.duty_cycle13(50),
		.output_clock_frequency14("0 MHz"),
		.phase_shift14("0 ps"),
		.duty_cycle14(50),
		.output_clock_frequency15("0 MHz"),
		.phase_shift15("0 ps"),
		.duty_cycle15(50),
		.output_clock_frequency16("0 MHz"),
		.phase_shift16("0 ps"),
		.duty_cycle16(50),
		.output_clock_frequency17("0 MHz"),
		.phase_shift17("0 ps"),
		.duty_cycle17(50),
		.pll_type("General"),
		.pll_subtype("General")
	) altera_pll_i (
		.rst	(areset),
		.outclk_0	(tx_hash_clk[0]),
		.outclk_1	(tx_hash_clk[1]),
		.locked	(lock),
		.fboutclk	( ),
		.fbclk	(1'b0),
		.refclk	(rx_clk)
	);

//	altpll	altpll_component (
//		.inclk ({1'b0, rx_clk}),
//		.clk (clks),
//		.activeclock (),
//		.areset (areset),
//		.clkbad (),
//		.clkena ({6{1'b1}}),
//		.clkloss (),
//		.clkswitch (1'b0),
//		.configupdate (1'b0),
//		.enable0 (),
//		.enable1 (),
//		.extclk (),
//		.extclkena ({4{1'b1}}),
//		.fbin (1'b1),
//		.fbmimicbidir (),
//		.fbout (),
//		.fref (),
//		.icdrclk (),
//		.locked (lock),
//		.pfdena (1'b1),
//		.phasecounterselect ({4{1'b1}}),
//		.phasedone (),
//		.phasestep (1'b1),
//		.phaseupdown (1'b1),
//		.pllena (1'b1),
//		.scanaclr (1'b0),
//		.scanclk (1'b0),
//		.scanclkena (1'b1),
//		.scandata (1'b0),
//		.scandataout (),
//		.scandone (),
//		.scanread (1'b0),
//		.scanwrite (1'b0),
//		.sclkout0 (),
//		.sclkout1 (),
//		.vcooverrange (),
//		.vcounderrange ());
//	defparam
//		altpll_component.bandwidth_type = "AUTO",
//		altpll_component.clk0_divide_by = DIVIDE_BY,
//		altpll_component.clk0_duty_cycle = 50,
//		altpll_component.clk0_multiply_by = MULTIPLY_BY,
//		altpll_component.clk0_phase_shift = "0",
//		altpll_component.compensate_clock = "CLK0",
//		altpll_component.inclk0_input_frequency = (1000000 / INPUT_FREQUENCY),
//		altpll_component.intended_device_family = "Cyclone V",
//		altpll_component.lpm_hint = "CBX_MODULE_PREFIX=main_pll",
//		altpll_component.lpm_type = "altpll",
//		altpll_component.operation_mode = "NORMAL",
//		altpll_component.pll_type = "AUTO",
//		altpll_component.port_activeclock = "PORT_UNUSED",
//		altpll_component.port_areset = "PORT_UNUSED",
//		altpll_component.port_clkbad0 = "PORT_UNUSED",
//		altpll_component.port_clkbad1 = "PORT_UNUSED",
//		altpll_component.port_clkloss = "PORT_UNUSED",
//		altpll_component.port_clkswitch = "PORT_UNUSED",
//		altpll_component.port_configupdate = "PORT_UNUSED",
//		altpll_component.port_fbin = "PORT_UNUSED",
//		altpll_component.port_inclk0 = "PORT_USED",
//		altpll_component.port_inclk1 = "PORT_UNUSED",
//		altpll_component.port_locked = "PORT_UNUSED",
//		altpll_component.port_pfdena = "PORT_UNUSED",
//		altpll_component.port_phasecounterselect = "PORT_UNUSED",
//		altpll_component.port_phasedone = "PORT_UNUSED",
//		altpll_component.port_phasestep = "PORT_UNUSED",
//		altpll_component.port_phaseupdown = "PORT_UNUSED",
//		altpll_component.port_pllena = "PORT_UNUSED",
//		altpll_component.port_scanaclr = "PORT_UNUSED",
//		altpll_component.port_scanclk = "PORT_UNUSED",
//		altpll_component.port_scanclkena = "PORT_UNUSED",
//		altpll_component.port_scandata = "PORT_UNUSED",
//		altpll_component.port_scandataout = "PORT_UNUSED",
//		altpll_component.port_scandone = "PORT_UNUSED",
//		altpll_component.port_scanread = "PORT_UNUSED",
//		altpll_component.port_scanwrite = "PORT_UNUSED",
//		altpll_component.port_clk0 = "PORT_USED",
//		altpll_component.port_clk1 = "PORT_UNUSED",
//		altpll_component.port_clk2 = "PORT_UNUSED",
//		altpll_component.port_clk3 = "PORT_UNUSED",
//		altpll_component.port_clk4 = "PORT_UNUSED",
//		altpll_component.port_clk5 = "PORT_UNUSED",
//		altpll_component.port_clkena0 = "PORT_UNUSED",
//		altpll_component.port_clkena1 = "PORT_UNUSED",
//		altpll_component.port_clkena2 = "PORT_UNUSED",
//		altpll_component.port_clkena3 = "PORT_UNUSED",
//		altpll_component.port_clkena4 = "PORT_UNUSED",
//		altpll_component.port_clkena5 = "PORT_UNUSED",
//		altpll_component.port_extclk0 = "PORT_UNUSED",
//		altpll_component.port_extclk1 = "PORT_UNUSED",
//		altpll_component.port_extclk2 = "PORT_UNUSED",
//		altpll_component.port_extclk3 = "PORT_UNUSED",
//		altpll_component.width_clock = 5;

endmodule

